//plug pmod-led on PMOD2 and pmod-switch on PMOD3

module switch( output LED );
      
  assign LED = 0;

endmodule
